module fpmul();
endmodule
