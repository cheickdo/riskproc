module fdiv(
    input clk,
    input resetn,
    input [31:0] rs1,
    input [31:0] rs2,
    output [31:0] out
);

wire [31:0] reciprocal;
endmodule