module fpcvt_from_int();
endmodule