module fpcvt_to_int();

endmodule