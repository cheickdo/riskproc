

module proc();

    //define internal processor bus here

    control c();
    datapath d();
endmodule
