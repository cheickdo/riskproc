module fpsqrt();
endmodule