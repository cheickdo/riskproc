module interrupt_ctrl();
endmodule