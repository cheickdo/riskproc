module csr(
    input clk,
    input [11:0] csr_addr
);
    reg [11:0] csreg [11:0];

endmodule