module dispatcher();
endmodule
