module fpaddsub();
endmodule