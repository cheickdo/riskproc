

module proc();
endmodule
