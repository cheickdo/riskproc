module fpdiv();
endmodule